module top;
    
endmodule